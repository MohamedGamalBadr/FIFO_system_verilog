package shared_pkg;
		logic test_finished;
		 int error_count = 0 , correct_count = 0 ;
	
endpackage